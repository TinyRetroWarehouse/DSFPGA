library ieee;
use ieee.std_logic_1164.all;

entity SyncRamDualByteEnable is
   generic 
   (
      BYTE_WIDTH : natural := 8;
      ADDR_WIDTH : natural := 6;
      BYTES      : natural := 4
   );
   port 
   (
      clk        : in std_logic;
      
      addr_a     : in natural range 0 to 2**ADDR_WIDTH - 1;
      datain_a0  : in std_logic_vector((BYTE_WIDTH-1) downto 0);
      datain_a1  : in std_logic_vector((BYTE_WIDTH-1) downto 0);
      datain_a2  : in std_logic_vector((BYTE_WIDTH-1) downto 0);
      datain_a3  : in std_logic_vector((BYTE_WIDTH-1) downto 0);
      dataout_a  : out std_logic_vector((BYTES*BYTE_WIDTH-1) downto 0) := (others => '0');
      we_a       : in std_logic := '1';
      be_a       : in  std_logic_vector (BYTES - 1 downto 0);
		            
      addr_b     : in natural range 0 to 2**ADDR_WIDTH - 1;
      datain_b0  : in std_logic_vector((BYTE_WIDTH-1) downto 0);
      datain_b1  : in std_logic_vector((BYTE_WIDTH-1) downto 0);
      datain_b2  : in std_logic_vector((BYTE_WIDTH-1) downto 0);
      datain_b3  : in std_logic_vector((BYTE_WIDTH-1) downto 0);
      dataout_b  : out std_logic_vector((BYTES*BYTE_WIDTH-1) downto 0) := (others => '0');
      we_b       : in std_logic := '1';
      be_b       : in  std_logic_vector (BYTES - 1 downto 0)
   );
end;

architecture rtl of SyncRamDualByteEnable is

	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(31 downto 0);
	signal ram : ram_t := (others => (others => '0'));
   
   signal addr_a_1 : natural range 0 to 2**ADDR_WIDTH - 1;
   signal addr_b_1 : natural range 0 to 2**ADDR_WIDTH - 1;
   signal we_a_1   : std_logic;
   signal we_b_1   : std_logic;

begin 
        
   process(clk)
   begin
      if(rising_edge(clk)) then 
      
         addr_a_1 <= addr_a;
         addr_b_1 <= addr_b;
         we_a_1   <= we_a;  
         we_b_1   <= we_b;  
      
         if(we_a = '1') then
            -- edit this code if using other than four bytes per word
            if(be_a(0) = '1') then
               ram(addr_a)(7 downto 0) <= datain_a0;
            end if;
            if be_a(1) = '1' then
               ram(addr_a)(15 downto 8) <= datain_a1;
            end if;
            if be_a(2) = '1' then
               ram(addr_a)(23 downto 16) <= datain_a2;
            end if;
            if be_a(3) = '1' then
               ram(addr_a)(31 downto 24) <= datain_a3;
            end if;
         end if;
         
         if (addr_a_1 /= addr_a or we_a_1 = '1' or we_b_1 = '1') then -- performance optimization for modelsim
            dataout_a <= ram(addr_a);
         end if;

         if(we_b = '1') then
               -- edit this code if using other than four bytes per word
            if(be_b(0) = '1') then
               ram(addr_b)(7 downto 0) <= datain_b0;
            end if;
            if be_b(1) = '1' then
               ram(addr_b)(15 downto 8) <= datain_b1;
            end if;
            if be_b(2) = '1' then
               ram(addr_b)(23 downto 16) <= datain_b2;
            end if;
            if be_b(3) = '1' then
               ram(addr_b)(31 downto 24) <= datain_b3;
            end if;
         end if;
         
         if (addr_b_1 /= addr_b or we_a_1 = '1' or we_b_1 = '1') then
            dataout_b <= ram(addr_b);
         end if;
         
         
      end if;
   end process;  
   
  
end rtl;